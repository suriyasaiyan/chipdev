module i_afifo#(
  parameter DATA_WIDTH = 32,
  parameter ADDR_WIDTH =  8
  )(
  input wclk, rclk
);
  
endmodule
